<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-21.0896,-4.16665,91.0104,-62.9748</PageViewport>
<gate>
<ID>2</ID>
<type>BE_DECODER_3x8</type>
<position>17.5,-21.5</position>
<input>
<ID>ENABLE</ID>7 </input>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>4 </input>
<output>
<ID>OUT_1</ID>21 </output>
<output>
<ID>OUT_2</ID>22 </output>
<output>
<ID>OUT_3</ID>27 </output>
<output>
<ID>OUT_4</ID>26 </output>
<output>
<ID>OUT_6</ID>20 </output>
<output>
<ID>OUT_7</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>34,-11</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>34,-13.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>34,-16</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>DE_TO</type>
<position>38,-16</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>14</ID>
<type>DE_TO</type>
<position>38,-11</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>16</ID>
<type>DE_TO</type>
<position>38,-13.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>9.5,-20</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>34.5,-33</position>
<input>
<ID>N_in0</ID>28 </input>
<input>
<ID>N_in1</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>DA_FROM</type>
<position>9.5,-22.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>22</ID>
<type>DA_FROM</type>
<position>9.5,-25</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>23</ID>
<type>AE_OR3</type>
<position>28.5,-33</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>26 </input>
<input>
<ID>IN_2</ID>27 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>24</ID>
<type>EE_VDD</type>
<position>10,-14</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_OR4</type>
<position>28.5,-21</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<input>
<ID>IN_2</ID>22 </input>
<input>
<ID>IN_3</ID>21 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>28</ID>
<type>DE_TO</type>
<position>39.5,-21</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F(x1,x2,x3)=Sm(1,2,6,7)</lparam></gate>
<gate>
<ID>30</ID>
<type>DE_TO</type>
<position>38.5,-33</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID G(x1,x2,x3)=Sm(3,4,7)</lparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>35,-21</position>
<input>
<ID>N_in0</ID>23 </input>
<input>
<ID>N_in1</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-11,36,-11</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-11,36,-11</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-13.5,36,-13.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-13.5,36,-13.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-16,36,-16</points>
<intersection>-16 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-16,36,-16</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36,-16,36,-16</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-20,14.5,-20</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>14.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>14.5,-23,14.5,-20</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-24,13,-22.5</points>
<intersection>-24 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-24,14.5,-24</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-22.5,13,-22.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-25,14.5,-25</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>14.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>14.5,-25,14.5,-25</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-25 1</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-18,10,-15</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-18,14.5,-18</points>
<connection>
<GID>2</GID>
<name>ENABLE</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-18,25.5,-18</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>OUT_7</name></connection>
<intersection>25.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25.5,-31,25.5,-18</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-18 1</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-20,23,-19</points>
<intersection>-20 1</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-20,25.5,-20</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20.5,-19,23,-19</points>
<connection>
<GID>2</GID>
<name>OUT_6</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-24,25.5,-24</points>
<connection>
<GID>26</GID>
<name>IN_3</name></connection>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-23,23,-22</points>
<intersection>-23 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-22,25.5,-22</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20.5,-23,23,-23</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32.5,-21,34,-21</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<connection>
<GID>36</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-33,23,-21</points>
<intersection>-33 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-21,23,-21</points>
<connection>
<GID>2</GID>
<name>OUT_4</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-33,25.5,-33</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-35,23,-22</points>
<intersection>-35 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-22,23,-22</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-35,25.5,-35</points>
<connection>
<GID>23</GID>
<name>IN_2</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-33,33.5,-33</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<connection>
<GID>19</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>36,-21,37.5,-21</points>
<connection>
<GID>36</GID>
<name>N_in1</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>35.5,-33,36.5,-33</points>
<connection>
<GID>19</GID>
<name>N_in1</name></connection>
<connection>
<GID>30</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,13.6541,112.1,-45.1541</PageViewport></page 1>
<page 2>
<PageViewport>0,13.6541,112.1,-45.1541</PageViewport></page 2>
<page 3>
<PageViewport>0,13.6541,112.1,-45.1541</PageViewport></page 3>
<page 4>
<PageViewport>0,13.6541,112.1,-45.1541</PageViewport></page 4>
<page 5>
<PageViewport>0,13.6541,112.1,-45.1541</PageViewport></page 5>
<page 6>
<PageViewport>0,13.6541,112.1,-45.1541</PageViewport></page 6>
<page 7>
<PageViewport>0,13.6541,112.1,-45.1541</PageViewport></page 7>
<page 8>
<PageViewport>0,13.6541,112.1,-45.1541</PageViewport></page 8>
<page 9>
<PageViewport>0,13.6541,112.1,-45.1541</PageViewport></page 9></circuit>