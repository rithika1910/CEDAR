<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-274.838,35.5026,-151.852,-29.0164</PageViewport>
<gate>
<ID>2</ID>
<type>GA_LED</type>
<position>-209.5,14</position>
<input>
<ID>N_in0</ID>5 </input>
<input>
<ID>N_in1</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AE_SMALL_INVERTER</type>
<position>-237.5,19.5</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_SMALL_INVERTER</type>
<position>-237.5,15</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND3</type>
<position>-227,18</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>6 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>16</ID>
<type>DA_FROM</type>
<position>-235,11.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>-247,15</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>-223,-0.5</position>
<gparam>LABEL_TEXT F(A,B,C,D)=A'B'C+ABD'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>DA_FROM</type>
<position>-246.5,19.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND3</type>
<position>-227,7</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>4 </input>
<input>
<ID>IN_2</ID>9 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>-246,5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_SMALL_INVERTER</type>
<position>-239,5</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AE_OR2</type>
<position>-215,13.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>-212.5,27</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>-212.5,24.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>-212.5,21.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>-212.5,18.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>-203.5,24.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>-203.5,18.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>-203.5,21.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>48</ID>
<type>DE_TO</type>
<position>-203.5,27</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>54</ID>
<type>DE_TO</type>
<position>-205,14</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F(A,B,C,D)</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-232.5,19.5,-232.5,20</points>
<intersection>19.5 2</intersection>
<intersection>20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-232.5,20,-230,20</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-232.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-235.5,19.5,-232.5,19.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-232.5,15,-232.5,18</points>
<intersection>15 2</intersection>
<intersection>18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-232.5,18,-230,18</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>-232.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-235.5,15,-232.5,15</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-245,15,-239.5,15</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-241 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-241,7,-241,15</points>
<intersection>7 5</intersection>
<intersection>15 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-241,7,-230,7</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-241 4</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-211,13.5,-211,14</points>
<intersection>13.5 1</intersection>
<intersection>14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-212,13.5,-211,13.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>-211 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-211,14,-210.5,14</points>
<connection>
<GID>2</GID>
<name>N_in0</name></connection>
<intersection>-211 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-231.5,11.5,-231.5,16</points>
<intersection>11.5 3</intersection>
<intersection>16 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-233,11.5,-231.5,11.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-231.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-231.5,16,-230,16</points>
<connection>
<GID>10</GID>
<name>IN_2</name></connection>
<intersection>-231.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-244.5,19.5,-239.5,19.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-242.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-242.5,9,-242.5,19.5</points>
<intersection>9 4</intersection>
<intersection>19.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-242.5,9,-230,9</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-242.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-244,5,-241,5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-237,5,-230,5</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-221,14.5,-221,18</points>
<intersection>14.5 1</intersection>
<intersection>18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-221,14.5,-218,14.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-221 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-224,18,-221,18</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>-221 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-221,7,-221,12.5</points>
<intersection>7 2</intersection>
<intersection>12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-221,12.5,-218,12.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>-221 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-224,7,-221,7</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>-221 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-208.5,14,-207,14</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-210.5,27,-205.5,27</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<connection>
<GID>48</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-210.5,24.5,-205.5,24.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<connection>
<GID>42</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-210.5,21.5,-205.5,21.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-210.5,18.5,-205.5,18.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,130.447,627.187,-198.578</PageViewport></page 1>
<page 2>
<PageViewport>0,130.447,627.187,-198.578</PageViewport></page 2>
<page 3>
<PageViewport>0,130.447,627.187,-198.578</PageViewport></page 3>
<page 4>
<PageViewport>0,130.447,627.187,-198.578</PageViewport></page 4>
<page 5>
<PageViewport>0,130.447,627.187,-198.578</PageViewport></page 5>
<page 6>
<PageViewport>0,130.447,627.187,-198.578</PageViewport></page 6>
<page 7>
<PageViewport>0,130.447,627.187,-198.578</PageViewport></page 7>
<page 8>
<PageViewport>0,130.447,627.187,-198.578</PageViewport></page 8>
<page 9>
<PageViewport>0,130.447,627.187,-198.578</PageViewport></page 9></circuit>