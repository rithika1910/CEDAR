<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-312.995,36.4681,-150.455,-14.8301</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND3</type>
<position>-237,21.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>6 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND3</type>
<position>-237,12</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>7 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND3</type>
<position>-236.5,2.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>7 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_OR3</type>
<position>-213.5,12</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>3 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>-241.5,-5</position>
<gparam>LABEL_TEXT F(A,B,C,D)=ABC+BCD+ACD</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>DA_FROM</type>
<position>-267,23.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>22</ID>
<type>DA_FROM</type>
<position>-267.5,17</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>-268,8</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>26</ID>
<type>DA_FROM</type>
<position>-268,3</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>-207,12</position>
<input>
<ID>N_in0</ID>8 </input>
<input>
<ID>N_in2</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>-215.5,31.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>-215.5,28.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>-215.5,25.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>-215.5,22.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>38</ID>
<type>DE_TO</type>
<position>-210.5,31.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>-210.5,28.5</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>-210.5,25.5</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>-210.5,22.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>-202.5,12</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F(A,B,C,D)</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-225.5,14,-225.5,21.5</points>
<intersection>14 1</intersection>
<intersection>21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-225.5,14,-216.5,14</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-225.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-234,21.5,-225.5,21.5</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>-225.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-234,12,-216.5,12</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<connection>
<GID>16</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-225,2.5,-225,10</points>
<intersection>2.5 2</intersection>
<intersection>10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-225,10,-216.5,10</points>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<intersection>-225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-233.5,2.5,-225,2.5</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>-225 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-265,23.5,-240,23.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-259 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-259,4.5,-259,23.5</points>
<intersection>4.5 3</intersection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-259,4.5,-239.5,4.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-259 2</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-250.5,17,-250.5,21.5</points>
<intersection>17 2</intersection>
<intersection>21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-250.5,21.5,-240,21.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-250.5 0</intersection>
<intersection>-246 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-265.5,17,-250.5,17</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-250.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-246,14,-246,21.5</points>
<intersection>14 4</intersection>
<intersection>21.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-246,14,-240,14</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-246 3</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-249,8,-249,19.5</points>
<intersection>8 2</intersection>
<intersection>19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-249,19.5,-240,19.5</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>-249 0</intersection>
<intersection>-247.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-266,8,-249,8</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-249 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-247.5,12,-247.5,19.5</points>
<intersection>12 4</intersection>
<intersection>19.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-247.5,12,-240,12</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-247.5 3</intersection>
<intersection>-245 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-245,2.5,-245,12</points>
<intersection>2.5 6</intersection>
<intersection>12 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-245,2.5,-239.5,2.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-245 5</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-247.5,0.5,-247.5,10</points>
<intersection>0.5 3</intersection>
<intersection>3 4</intersection>
<intersection>10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-247.5,10,-240,10</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<intersection>-247.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-247.5,0.5,-239.5,0.5</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<intersection>-247.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-266,3,-247.5,3</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-247.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-210.5,12,-208,12</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<connection>
<GID>28</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-213.5,31.5,-212.5,31.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-213.5,28.5,-212.5,28.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-212.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-212.5,28.5,-212.5,28.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>28.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-213.5,25.5,-212.5,25.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>-212.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-212.5,25.5,-212.5,25.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>25.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-213.5,22.5,-212.5,22.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>-212.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-212.5,22.5,-212.5,22.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-207,11,-207,12</points>
<connection>
<GID>28</GID>
<name>N_in2</name></connection>
<intersection>12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-207,12,-204.5,12</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>-207 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,130.447,621.676,-65.7554</PageViewport></page 1>
<page 2>
<PageViewport>0,130.447,621.676,-65.7554</PageViewport></page 2>
<page 3>
<PageViewport>0,130.447,621.676,-65.7554</PageViewport></page 3>
<page 4>
<PageViewport>0,130.447,621.676,-65.7554</PageViewport></page 4>
<page 5>
<PageViewport>0,130.447,621.676,-65.7554</PageViewport></page 5>
<page 6>
<PageViewport>0,130.447,621.676,-65.7554</PageViewport></page 6>
<page 7>
<PageViewport>0,130.447,621.676,-65.7554</PageViewport></page 7>
<page 8>
<PageViewport>0,130.447,621.676,-65.7554</PageViewport></page 8>
<page 9>
<PageViewport>0,130.447,621.676,-65.7554</PageViewport></page 9></circuit>