<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-51.75,2.4167,62.05,-57.2833</PageViewport>
<gate>
<ID>194</ID>
<type>AA_LABEL</type>
<position>-29,-13</position>
<gparam>LABEL_TEXT y0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>197</ID>
<type>AA_LABEL</type>
<position>-29,-24.5</position>
<gparam>LABEL_TEXT y1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>199</ID>
<type>AA_LABEL</type>
<position>2.5,-36</position>
<gparam>LABEL_TEXT circuit for driving display</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>-42.5,-2</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>-42.5,-4.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>-42.5,-9.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>-42.5,-7</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>DE_TO</type>
<position>-36.5,-4.5</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID milk</lparam></gate>
<gate>
<ID>18</ID>
<type>DE_TO</type>
<position>-36.5,-7</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID tea</lparam></gate>
<gate>
<ID>20</ID>
<type>DE_TO</type>
<position>-36.5,-9.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID coffee</lparam></gate>
<gate>
<ID>22</ID>
<type>DE_TO</type>
<position>-36.5,-2</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cocoa</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>-41.5,-13.5</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID tea</lparam></gate>
<gate>
<ID>26</ID>
<type>DA_FROM</type>
<position>-41.5,-19.5</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cocoa</lparam></gate>
<gate>
<ID>28</ID>
<type>DA_FROM</type>
<position>-42,-27</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID milk</lparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>52,-11</position>
<input>
<ID>N_in1</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>54,-11</position>
<input>
<ID>N_in0</ID>15 </input>
<input>
<ID>N_in1</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>GA_LED</type>
<position>56,-11</position>
<input>
<ID>N_in0</ID>14 </input>
<input>
<ID>N_in1</ID>94 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>GA_LED</type>
<position>50,-13</position>
<input>
<ID>N_in2</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>GA_LED</type>
<position>50,-15</position>
<input>
<ID>N_in2</ID>16 </input>
<input>
<ID>N_in3</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>GA_LED</type>
<position>52,-19</position>
<input>
<ID>N_in0</ID>113 </input>
<input>
<ID>N_in1</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>GA_LED</type>
<position>58,-15</position>
<input>
<ID>N_in2</ID>11 </input>
<input>
<ID>N_in3</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>58,-13</position>
<input>
<ID>N_in2</ID>13 </input>
<input>
<ID>N_in3</ID>105 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>GA_LED</type>
<position>58,-17</position>
<input>
<ID>N_in2</ID>104 </input>
<input>
<ID>N_in3</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>GA_LED</type>
<position>56,-19</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>GA_LED</type>
<position>54,-19</position>
<input>
<ID>N_in0</ID>10 </input>
<input>
<ID>N_in1</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>GA_LED</type>
<position>50,-17</position>
<input>
<ID>N_in2</ID>99 </input>
<input>
<ID>N_in3</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>GA_LED</type>
<position>50,-21</position>
<input>
<ID>N_in0</ID>119 </input>
<input>
<ID>N_in2</ID>25 </input>
<input>
<ID>N_in3</ID>99 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>GA_LED</type>
<position>50,-23</position>
<input>
<ID>N_in2</ID>24 </input>
<input>
<ID>N_in3</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>GA_LED</type>
<position>52,-27</position>
<input>
<ID>N_in0</ID>101 </input>
<input>
<ID>N_in1</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>GA_LED</type>
<position>58,-23</position>
<input>
<ID>N_in2</ID>26 </input>
<input>
<ID>N_in3</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>GA_LED</type>
<position>58,-21</position>
<input>
<ID>N_in2</ID>27 </input>
<input>
<ID>N_in3</ID>104 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>GA_LED</type>
<position>58,-25</position>
<input>
<ID>N_in3</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>GA_LED</type>
<position>56,-27</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>GA_LED</type>
<position>54,-27</position>
<input>
<ID>N_in0</ID>19 </input>
<input>
<ID>N_in1</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>GA_LED</type>
<position>50,-25</position>
<input>
<ID>N_in3</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AO_XNOR2</type>
<position>3.5,-10</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>AE_OR2</type>
<position>-34.5,-14.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>AE_OR2</type>
<position>-34.5,-26</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>87</ID>
<type>AA_AND2</type>
<position>3.5,-15.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>AI_XOR2</type>
<position>4,-32</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>91</ID>
<type>AE_OR2</type>
<position>14.5,-26</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_AND2</type>
<position>4,-25</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>97</ID>
<type>AE_SMALL_INVERTER</type>
<position>-10,-26</position>
<input>
<ID>IN_0</ID>37 </input>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>99</ID>
<type>AE_SMALL_INVERTER</type>
<position>-10,-24</position>
<input>
<ID>IN_0</ID>38 </input>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>103</ID>
<type>AE_OR2</type>
<position>14.5,-20</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>105</ID>
<type>AE_OR2</type>
<position>14,-3.5</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_AND2</type>
<position>3.5,-2.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>130</ID>
<type>DA_FROM</type>
<position>-41.5,-33.5</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID tea</lparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>-41.5,-37.5</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID cocoa</lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>-41.5,-35.5</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID milk</lparam></gate>
<gate>
<ID>135</ID>
<type>DA_FROM</type>
<position>-41.5,-31.5</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID coffee</lparam></gate>
<gate>
<ID>147</ID>
<type>AM_MUX_16x1</type>
<position>-28.5,-48</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>89 </input>
<input>
<ID>IN_10</ID>90 </input>
<input>
<ID>IN_11</ID>90 </input>
<input>
<ID>IN_12</ID>90 </input>
<input>
<ID>IN_13</ID>90 </input>
<input>
<ID>IN_14</ID>90 </input>
<input>
<ID>IN_15</ID>90 </input>
<input>
<ID>IN_2</ID>89 </input>
<input>
<ID>IN_3</ID>90 </input>
<input>
<ID>IN_4</ID>89 </input>
<input>
<ID>IN_5</ID>90 </input>
<input>
<ID>IN_6</ID>90 </input>
<input>
<ID>IN_7</ID>90 </input>
<input>
<ID>IN_8</ID>89 </input>
<input>
<ID>IN_9</ID>90 </input>
<output>
<ID>OUT</ID>93 </output>
<input>
<ID>SEL_0</ID>83 </input>
<input>
<ID>SEL_1</ID>84 </input>
<input>
<ID>SEL_2</ID>87 </input>
<input>
<ID>SEL_3</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>149</ID>
<type>EE_VDD</type>
<position>-48.5,-42</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>153</ID>
<type>FF_GND</type>
<position>-43,-46</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_AND2</type>
<position>34.5,-11</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_AND2</type>
<position>34.5,-16.5</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_AND2</type>
<position>34.5,-21</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_AND2</type>
<position>34.5,-27</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>165</ID>
<type>AA_AND2</type>
<position>34.5,-4.5</position>
<input>
<ID>IN_0</ID>114 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_LABEL</type>
<position>53.5,-9</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_LABEL</type>
<position>38,-10</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>AA_LABEL</type>
<position>60,-15</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AA_LABEL</type>
<position>60,-22.5</position>
<gparam>LABEL_TEXT c</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>AA_LABEL</type>
<position>54.5,-29</position>
<gparam>LABEL_TEXT d</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>AA_LABEL</type>
<position>48,-22.5</position>
<gparam>LABEL_TEXT e</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>AA_LABEL</type>
<position>48,-15</position>
<gparam>LABEL_TEXT f</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>AA_LABEL</type>
<position>54,-20.5</position>
<gparam>LABEL_TEXT g</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_LABEL</type>
<position>39,-15.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>40.5,-15.5</position>
<gparam>LABEL_TEXT c</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>AA_LABEL</type>
<position>38.5,-3</position>
<gparam>LABEL_TEXT g</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>38.5,-26</position>
<gparam>LABEL_TEXT d</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>AA_LABEL</type>
<position>39,-20</position>
<gparam>LABEL_TEXT e</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>188</ID>
<type>AA_LABEL</type>
<position>40.5,-20</position>
<gparam>LABEL_TEXT f</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>AA_LABEL</type>
<position>-35.5,-29</position>
<gparam>LABEL_TEXT Encoder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>192</ID>
<type>AA_LABEL</type>
<position>-24.5,-47</position>
<gparam>LABEL_TEXT f</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40.5,-2,-38.5,-2</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<connection>
<GID>22</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40.5,-4.5,-38.5,-4.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<connection>
<GID>16</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40.5,-7,-38.5,-7</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40.5,-9.5,-38.5,-9.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>55,-19,55,-19</points>
<connection>
<GID>50</GID>
<name>N_in0</name></connection>
<connection>
<GID>51</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>53,-19,53,-19</points>
<connection>
<GID>46</GID>
<name>N_in1</name></connection>
<connection>
<GID>51</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-16,58,-16</points>
<connection>
<GID>47</GID>
<name>N_in2</name></connection>
<connection>
<GID>49</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-14,58,-14</points>
<connection>
<GID>47</GID>
<name>N_in3</name></connection>
<connection>
<GID>48</GID>
<name>N_in2</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-11,55,-11</points>
<connection>
<GID>38</GID>
<name>N_in1</name></connection>
<connection>
<GID>40</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-11,53,-11</points>
<connection>
<GID>36</GID>
<name>N_in1</name></connection>
<connection>
<GID>38</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>50,-16,50,-16</points>
<connection>
<GID>44</GID>
<name>N_in2</name></connection>
<connection>
<GID>57</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>50,-14,50,-14</points>
<connection>
<GID>42</GID>
<name>N_in2</name></connection>
<connection>
<GID>44</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>55,-27,55,-27</points>
<connection>
<GID>71</GID>
<name>N_in0</name></connection>
<connection>
<GID>72</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>53,-27,53,-27</points>
<connection>
<GID>67</GID>
<name>N_in1</name></connection>
<connection>
<GID>72</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>50,-24,50,-24</points>
<connection>
<GID>66</GID>
<name>N_in2</name></connection>
<connection>
<GID>73</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>50,-22,50,-22</points>
<connection>
<GID>65</GID>
<name>N_in2</name></connection>
<connection>
<GID>66</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-24,58,-24</points>
<connection>
<GID>68</GID>
<name>N_in2</name></connection>
<connection>
<GID>70</GID>
<name>N_in3</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-22,58,-22</points>
<connection>
<GID>68</GID>
<name>N_in3</name></connection>
<connection>
<GID>69</GID>
<name>N_in2</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-39.5,-13.5,-37.5,-13.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<connection>
<GID>77</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-39.5,-19.5,-37.5,-19.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-37.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-37.5,-25,-37.5,-15.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>-19.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-27,-37.5,-27</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<connection>
<GID>79</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,-33,-19.5,-11</points>
<intersection>-33 6</intersection>
<intersection>-26 4</intersection>
<intersection>-16.5 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-19.5,-11,0.5,-11</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-16.5,0.5,-16.5</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-31.5,-26,-12,-26</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-19.5,-33,1,-33</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-9,0.5,-9</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>-6.5 2</intersection>
<intersection>-5.5 9</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-6.5,-14.5,-6.5,-9</points>
<intersection>-14.5 3</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-31.5,-14.5,0.5,-14.5</points>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>-13.5 4</intersection>
<intersection>-12 14</intersection>
<intersection>-6.5 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-13.5,-31,-13.5,-14.5</points>
<intersection>-31 8</intersection>
<intersection>-14.5 3</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-13.5,-31,1,-31</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>-13.5 4</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-5.5,-9,-5.5,-1.5</points>
<intersection>-9 1</intersection>
<intersection>-1.5 16</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-12,-24,-12,-14.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>-14.5 3</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-5.5,-1.5,0.5,-1.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>-5.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-32,8,-21</points>
<intersection>-32 5</intersection>
<intersection>-27 1</intersection>
<intersection>-21 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-27,11.5,-27</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>8,-21,11.5,-21</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>7,-32,8,-32</points>
<connection>
<GID>89</GID>
<name>OUT</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>7,-25,11.5,-25</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<connection>
<GID>95</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8,-24,1,-24</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8,-26,1,-26</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>-4 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-4,-26,-4,-3.5</points>
<intersection>-26 1</intersection>
<intersection>-3.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-4,-3.5,0.5,-3.5</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>-4 2</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27,-38.5,-27,-31.5</points>
<connection>
<GID>147</GID>
<name>SEL_0</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39.5,-31.5,-27,-31.5</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>-27 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-38.5,-28,-33.5</points>
<connection>
<GID>147</GID>
<name>SEL_1</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39.5,-33.5,-28,-33.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>-28 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-38.5,-30,-37.5</points>
<connection>
<GID>147</GID>
<name>SEL_3</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39.5,-37.5,-30,-37.5</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-38.5,-29,-35.5</points>
<connection>
<GID>147</GID>
<name>SEL_2</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39.5,-35.5,-29,-35.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48.5,-47.5,-48.5,-43</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,-47.5,-31.5,-47.5</points>
<connection>
<GID>147</GID>
<name>IN_8</name></connection>
<intersection>-48.5 0</intersection>
<intersection>-31.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-31.5,-54.5,-31.5,-47.5</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<connection>
<GID>147</GID>
<name>IN_2</name></connection>
<connection>
<GID>147</GID>
<name>IN_4</name></connection>
<intersection>-47.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-46.5,-43,-45</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-43,-46.5,-31.5,-46.5</points>
<connection>
<GID>147</GID>
<name>IN_9</name></connection>
<intersection>-43 0</intersection>
<intersection>-31.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-31.5,-55.5,-31.5,-40.5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<connection>
<GID>147</GID>
<name>IN_10</name></connection>
<connection>
<GID>147</GID>
<name>IN_11</name></connection>
<connection>
<GID>147</GID>
<name>IN_12</name></connection>
<connection>
<GID>147</GID>
<name>IN_13</name></connection>
<connection>
<GID>147</GID>
<name>IN_14</name></connection>
<connection>
<GID>147</GID>
<name>IN_3</name></connection>
<connection>
<GID>147</GID>
<name>IN_5</name></connection>
<connection>
<GID>147</GID>
<name>IN_6</name></connection>
<connection>
<GID>147</GID>
<name>IN_7</name></connection>
<connection>
<GID>147</GID>
<name>IN_15</name></connection>
<intersection>-46.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6.5,-10,8,-10</points>
<connection>
<GID>75</GID>
<name>OUT</name></connection>
<intersection>8 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>8,-19,8,-10</points>
<intersection>-19 4</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>8,-19,31.5,-19</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>8 3</intersection>
<intersection>31.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>31.5,-26,31.5,-19</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>-19 4</intersection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-22,27.5,-5.5</points>
<intersection>-22 8</intersection>
<intersection>-17.5 3</intersection>
<intersection>-12 11</intersection>
<intersection>-5.5 12</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-25.5,-17.5,27.5,-17.5</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>-25.5 13</intersection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>27.5,-22,31.5,-22</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection>
<intersection>31.5 14</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>27.5,-12,31.5,-12</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>27.5,-5.5,31.5,-5.5</points>
<connection>
<GID>165</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-25.5,-48,-25.5,-17.5</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<intersection>-17.5 3</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>31.5,-28,31.5,-22</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<intersection>-22 8</intersection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>37.5,-11,57,-11</points>
<connection>
<GID>155</GID>
<name>OUT</name></connection>
<connection>
<GID>40</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>17.5,-20,31.5,-20</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<connection>
<GID>103</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-20,50,-18</points>
<connection>
<GID>57</GID>
<name>N_in2</name></connection>
<connection>
<GID>65</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>17.5,-26,31.5,-26</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<connection>
<GID>91</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>37.5,-27,51,-27</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<connection>
<GID>67</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6.5,-2.5,11,-2.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<connection>
<GID>107</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-15.5,10.5,-4.5</points>
<intersection>-15.5 1</intersection>
<intersection>-15.5 1</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-15.5,31.5,-15.5</points>
<connection>
<GID>87</GID>
<name>OUT</name></connection>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10.5,-4.5,11,-4.5</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-20,58,-18</points>
<connection>
<GID>49</GID>
<name>N_in2</name></connection>
<connection>
<GID>69</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-16.5,58,-12</points>
<connection>
<GID>48</GID>
<name>N_in3</name></connection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-16.5,58,-16.5</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-19,44,-4.5</points>
<intersection>-19 4</intersection>
<intersection>-4.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>37.5,-4.5,44,-4.5</points>
<connection>
<GID>165</GID>
<name>OUT</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>44,-19,51,-19</points>
<connection>
<GID>46</GID>
<name>N_in0</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>17,-3.5,31.5,-3.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<connection>
<GID>105</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>37.5,-21,49,-21</points>
<connection>
<GID>159</GID>
<name>OUT</name></connection>
<connection>
<GID>65</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,6.2852e-007,113.8,-59.7</PageViewport></page 1>
<page 2>
<PageViewport>0,6.2852e-007,113.8,-59.7</PageViewport></page 2>
<page 3>
<PageViewport>0,6.2852e-007,113.8,-59.7</PageViewport></page 3>
<page 4>
<PageViewport>0,6.2852e-007,113.8,-59.7</PageViewport></page 4>
<page 5>
<PageViewport>0,6.2852e-007,113.8,-59.7</PageViewport></page 5>
<page 6>
<PageViewport>0,6.2852e-007,113.8,-59.7</PageViewport></page 6>
<page 7>
<PageViewport>0,6.2852e-007,113.8,-59.7</PageViewport></page 7>
<page 8>
<PageViewport>0,6.2852e-007,113.8,-59.7</PageViewport></page 8>
<page 9>
<PageViewport>0,6.2852e-007,113.8,-59.7</PageViewport></page 9></circuit>