<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-11.7333,-5.1,101.667,-46.2</PageViewport>
<gate>
<ID>2</ID>
<type>AA_MUX_2x1</type>
<position>33,-15.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>1 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_MUX_4x1</type>
<position>46.5,-30</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_2</ID>13 </input>
<input>
<ID>IN_3</ID>1 </input>
<output>
<ID>OUT</ID>2 </output>
<input>
<ID>SEL_0</ID>23 </input>
<input>
<ID>SEL_1</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>53,-21.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>55,-30</position>
<input>
<ID>N_in0</ID>2 </input>
<input>
<ID>N_in1</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>53,-16.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>53,-19</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>53,-24</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>16</ID>
<type>EE_VDD</type>
<position>26.5,-13</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>18</ID>
<type>DE_TO</type>
<position>58.5,-16.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>20</ID>
<type>DE_TO</type>
<position>58.5,-19</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>22</ID>
<type>DE_TO</type>
<position>58.5,-21.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>24</ID>
<type>DE_TO</type>
<position>58.5,-24</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_SMALL_INVERTER</type>
<position>27.5,-16.5</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>28</ID>
<type>DA_FROM</type>
<position>21,-16.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>30.5,-33</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x4</lparam></gate>
<gate>
<ID>32</ID>
<type>DA_FROM</type>
<position>31,-29</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>34</ID>
<type>AE_SMALL_INVERTER</type>
<position>36.5,-31</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>31,-9.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x1</lparam></gate>
<gate>
<ID>38</ID>
<type>DA_FROM</type>
<position>44.5,-21</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x3</lparam></gate>
<gate>
<ID>40</ID>
<type>DA_FROM</type>
<position>44.5,-23.5</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID x2</lparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>58,-30</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID f(x1,x2,x3,x4)</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>45,-37</position>
<gparam>LABEL_TEXT f(x1,x2,x3,x4) = x2'x3'x4+x3x4'+x1x2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-27,39,-15.5</points>
<intersection>-27 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-27,43.5,-27</points>
<connection>
<GID>4</GID>
<name>IN_3</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-15.5,39,-15.5</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-30,54,-30</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<connection>
<GID>8</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-14.5,26.5,-14</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-14.5,31,-14.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-16.5,56.5,-16.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>56.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>56.5,-16.5,56.5,-16.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-16.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-19,56.5,-19</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-21.5,56.5,-21.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>22</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-24,56.5,-24</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-16.5,31,-16.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-16.5,25.5,-16.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32.5,-33,43.5,-33</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>34.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>34.5,-33,34.5,-31</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>-33 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-31,43.5,-31</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33,-29,43.5,-29</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>33,-13,33,-9.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-30,56,-30</points>
<connection>
<GID>8</GID>
<name>N_in1</name></connection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-30,56,-30</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-25,46.5,-23.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>SEL_1</name></connection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-25,47.5,-21</points>
<connection>
<GID>4</GID>
<name>SEL_0</name></connection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-21,47.5,-21</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,113.4,-41.1</PageViewport></page 1>
<page 2>
<PageViewport>0,0,113.4,-41.1</PageViewport></page 2>
<page 3>
<PageViewport>0,0,113.4,-41.1</PageViewport></page 3>
<page 4>
<PageViewport>0,0,113.4,-41.1</PageViewport></page 4>
<page 5>
<PageViewport>0,0,113.4,-41.1</PageViewport></page 5>
<page 6>
<PageViewport>0,0,113.4,-41.1</PageViewport></page 6>
<page 7>
<PageViewport>0,0,113.4,-41.1</PageViewport></page 7>
<page 8>
<PageViewport>0,0,113.4,-41.1</PageViewport></page 8>
<page 9>
<PageViewport>0,0,113.4,-41.1</PageViewport></page 9></circuit>