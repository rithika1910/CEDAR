<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-13.402,-3.40811,86.7629,-28.9802</PageViewport>
<gate>
<ID>2</ID>
<type>DE_TO</type>
<position>45.5,-20.5</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F(a,b,c,d)</lparam></gate>
<gate>
<ID>5</ID>
<type>BA_NAND2</type>
<position>24,-20.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>BA_NAND2</type>
<position>22.5,-15.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>BA_NAND3</type>
<position>36,-20.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>12 </input>
<input>
<ID>IN_2</ID>20 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>10</ID>
<type>DA_FROM</type>
<position>6.5,-14.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a</lparam></gate>
<gate>
<ID>11</ID>
<type>BA_NAND2</type>
<position>21,-25.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>DA_FROM</type>
<position>6.5,-21.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c</lparam></gate>
<gate>
<ID>14</ID>
<type>DA_FROM</type>
<position>6.5,-18</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b</lparam></gate>
<gate>
<ID>16</ID>
<type>DA_FROM</type>
<position>6.5,-24.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID d</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>54.5,-5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>54.5,-8</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>54.5,-11</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>54.5,-14</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>42.5,-20.5</position>
<input>
<ID>N_in0</ID>14 </input>
<input>
<ID>N_in1</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>61.5,-5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID a</lparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>61.5,-8</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID b</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>61.5,-11</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID c</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>61.5,-14</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID d</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-14.5,19.5,-14.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>16.5 7</intersection>
<intersection>19.5 9</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>16.5,-21.5,16.5,-14.5</points>
<intersection>-21.5 8</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>16.5,-21.5,21,-21.5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>16.5 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>19.5,-14.5,19.5,-14.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-21.5,14,-21.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>14 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>14,-21.5,14,-16.5</points>
<intersection>-21.5 1</intersection>
<intersection>-16.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>14,-16.5,19.5,-16.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>14 4</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>43.5,-20.5,43.5,-20.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>38</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-19.5,14.5,-18</points>
<intersection>-19.5 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-18,14.5,-18</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-19.5,21,-19.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-18.5,29,-15.5</points>
<intersection>-18.5 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-18.5,33,-18.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-15.5,29,-15.5</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-20.5,33,-20.5</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<connection>
<GID>8</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-20.5,41.5,-20.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<connection>
<GID>38</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-24.5,18,-24.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>18 3</intersection>
<intersection>18 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>18,-26.5,18,-24.5</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>18,-24.5,18,-24.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>-24.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56.5,-5,59.5,-5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>56.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>56.5,-5,56.5,-5</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>-5 1</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56.5,-8,59.5,-8</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>59.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>59.5,-8,59.5,-8</points>
<intersection>-8 1</intersection>
<intersection>-8 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59.5,-8,59.5,-8</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>59.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56.5,-11,59.5,-11</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>59.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>59.5,-11,59.5,-11</points>
<intersection>-11 1</intersection>
<intersection>-11 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>59.5,-11,59.5,-11</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>59.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56.5,-14,59.5,-14</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>59.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>59.5,-14,59.5,-14</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>-14 1</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-25.5,28.5,-22.5</points>
<intersection>-25.5 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-22.5,33,-22.5</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-25.5,28.5,-25.5</points>
<connection>
<GID>11</GID>
<name>OUT</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,105.438,750.388,-86.1364</PageViewport></page 1>
<page 2>
<PageViewport>0,105.438,750.388,-86.1364</PageViewport></page 2>
<page 3>
<PageViewport>0,105.438,750.388,-86.1364</PageViewport></page 3>
<page 4>
<PageViewport>0,105.438,750.388,-86.1364</PageViewport></page 4>
<page 5>
<PageViewport>0,105.438,750.388,-86.1364</PageViewport></page 5>
<page 6>
<PageViewport>0,105.438,750.388,-86.1364</PageViewport></page 6>
<page 7>
<PageViewport>0,105.438,750.388,-86.1364</PageViewport></page 7>
<page 8>
<PageViewport>0,105.438,750.388,-86.1364</PageViewport></page 8>
<page 9>
<PageViewport>0,105.438,750.388,-86.1364</PageViewport></page 9></circuit>